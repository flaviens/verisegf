module sub;
endmodule

module mid_a;
  sub i_sub;
endmodule

module sub;
endmodule

module mid_b;
  sub i_sub;
endmodule

module top;
  mid_a a;
  mid_b b;
endmodule
